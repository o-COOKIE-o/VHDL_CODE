--Last Update 2025.11.08 by COOKIE
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_arith.all;
use IEEE.std_logic_unsigned.all;

package typ is
  type slv1_vector   is array (natural range<>) of std_logic_vector(  0 downto 0);
  type slv2_vector   is array (natural range<>) of std_logic_vector(  1 downto 0);
  type slv3_vector   is array (natural range<>) of std_logic_vector(  2 downto 0);
  type slv4_vector   is array (natural range<>) of std_logic_vector(  3 downto 0);
  type slv5_vector   is array (natural range<>) of std_logic_vector(  4 downto 0);
  type slv6_vector   is array (natural range<>) of std_logic_vector(  5 downto 0);
  type slv7_vector   is array (natural range<>) of std_logic_vector(  6 downto 0);
  type slv8_vector   is array (natural range<>) of std_logic_vector(  7 downto 0);
  type slv9_vector   is array (natural range<>) of std_logic_vector(  8 downto 0);
  type slv10_vector  is array (natural range<>) of std_logic_vector(  9 downto 0);
  type slv11_vector  is array (natural range<>) of std_logic_vector( 10 downto 0);
  type slv12_vector  is array (natural range<>) of std_logic_vector( 11 downto 0);
  type slv13_vector  is array (natural range<>) of std_logic_vector( 12 downto 0);
  type slv14_vector  is array (natural range<>) of std_logic_vector( 13 downto 0);
  type slv15_vector  is array (natural range<>) of std_logic_vector( 14 downto 0);
  type slv16_vector  is array (natural range<>) of std_logic_vector( 15 downto 0);
  type slv17_vector  is array (natural range<>) of std_logic_vector( 16 downto 0);
  type slv18_vector  is array (natural range<>) of std_logic_vector( 17 downto 0);
  type slv19_vector  is array (natural range<>) of std_logic_vector( 18 downto 0);
  type slv20_vector  is array (natural range<>) of std_logic_vector( 19 downto 0);
  type slv21_vector  is array (natural range<>) of std_logic_vector( 20 downto 0);
  type slv22_vector  is array (natural range<>) of std_logic_vector( 21 downto 0);
  type slv23_vector  is array (natural range<>) of std_logic_vector( 22 downto 0);
  type slv24_vector  is array (natural range<>) of std_logic_vector( 23 downto 0);
  type slv25_vector  is array (natural range<>) of std_logic_vector( 24 downto 0);
  type slv26_vector  is array (natural range<>) of std_logic_vector( 25 downto 0);
  type slv27_vector  is array (natural range<>) of std_logic_vector( 26 downto 0);
  type slv28_vector  is array (natural range<>) of std_logic_vector( 27 downto 0);
  type slv29_vector  is array (natural range<>) of std_logic_vector( 28 downto 0);
  type slv30_vector  is array (natural range<>) of std_logic_vector( 29 downto 0);
  type slv31_vector  is array (natural range<>) of std_logic_vector( 30 downto 0);
  type slv32_vector  is array (natural range<>) of std_logic_vector( 31 downto 0);
  type slv33_vector  is array (natural range<>) of std_logic_vector( 32 downto 0);
  type slv34_vector  is array (natural range<>) of std_logic_vector( 33 downto 0);
  type slv35_vector  is array (natural range<>) of std_logic_vector( 34 downto 0);
  type slv36_vector  is array (natural range<>) of std_logic_vector( 35 downto 0);
  type slv37_vector  is array (natural range<>) of std_logic_vector( 36 downto 0);
  type slv38_vector  is array (natural range<>) of std_logic_vector( 37 downto 0);
  type slv39_vector  is array (natural range<>) of std_logic_vector( 38 downto 0);
  type slv40_vector  is array (natural range<>) of std_logic_vector( 39 downto 0);
  type slv41_vector  is array (natural range<>) of std_logic_vector( 40 downto 0);
  type slv42_vector  is array (natural range<>) of std_logic_vector( 41 downto 0);
  type slv43_vector  is array (natural range<>) of std_logic_vector( 42 downto 0);
  type slv44_vector  is array (natural range<>) of std_logic_vector( 43 downto 0);
  type slv45_vector  is array (natural range<>) of std_logic_vector( 44 downto 0);
  type slv46_vector  is array (natural range<>) of std_logic_vector( 45 downto 0);
  type slv47_vector  is array (natural range<>) of std_logic_vector( 46 downto 0);
  type slv48_vector  is array (natural range<>) of std_logic_vector( 47 downto 0);
  type slv49_vector  is array (natural range<>) of std_logic_vector( 48 downto 0);
  type slv50_vector  is array (natural range<>) of std_logic_vector( 49 downto 0);
  type slv51_vector  is array (natural range<>) of std_logic_vector( 50 downto 0);
  type slv52_vector  is array (natural range<>) of std_logic_vector( 51 downto 0);
  type slv53_vector  is array (natural range<>) of std_logic_vector( 52 downto 0);
  type slv54_vector  is array (natural range<>) of std_logic_vector( 53 downto 0);
  type slv55_vector  is array (natural range<>) of std_logic_vector( 54 downto 0);
  type slv56_vector  is array (natural range<>) of std_logic_vector( 55 downto 0);
  type slv57_vector  is array (natural range<>) of std_logic_vector( 56 downto 0);
  type slv58_vector  is array (natural range<>) of std_logic_vector( 57 downto 0);
  type slv59_vector  is array (natural range<>) of std_logic_vector( 58 downto 0);
  type slv60_vector  is array (natural range<>) of std_logic_vector( 59 downto 0);
  type slv61_vector  is array (natural range<>) of std_logic_vector( 60 downto 0);
  type slv62_vector  is array (natural range<>) of std_logic_vector( 61 downto 0);
  type slv63_vector  is array (natural range<>) of std_logic_vector( 62 downto 0);
  type slv64_vector  is array (natural range<>) of std_logic_vector( 63 downto 0);
  type slv65_vector  is array (natural range<>) of std_logic_vector( 64 downto 0);
  type slv66_vector  is array (natural range<>) of std_logic_vector( 65 downto 0);
  type slv67_vector  is array (natural range<>) of std_logic_vector( 66 downto 0);
  type slv68_vector  is array (natural range<>) of std_logic_vector( 67 downto 0);
  type slv69_vector  is array (natural range<>) of std_logic_vector( 68 downto 0);
  type slv70_vector  is array (natural range<>) of std_logic_vector( 69 downto 0);
  type slv71_vector  is array (natural range<>) of std_logic_vector( 70 downto 0);
  type slv72_vector  is array (natural range<>) of std_logic_vector( 71 downto 0);
  type slv73_vector  is array (natural range<>) of std_logic_vector( 72 downto 0);
  type slv74_vector  is array (natural range<>) of std_logic_vector( 73 downto 0);
  type slv75_vector  is array (natural range<>) of std_logic_vector( 74 downto 0);
  type slv76_vector  is array (natural range<>) of std_logic_vector( 75 downto 0);
  type slv77_vector  is array (natural range<>) of std_logic_vector( 76 downto 0);
  type slv78_vector  is array (natural range<>) of std_logic_vector( 77 downto 0);
  type slv79_vector  is array (natural range<>) of std_logic_vector( 78 downto 0);
  type slv80_vector  is array (natural range<>) of std_logic_vector( 79 downto 0);
  type slv81_vector  is array (natural range<>) of std_logic_vector( 80 downto 0);
  type slv82_vector  is array (natural range<>) of std_logic_vector( 81 downto 0);
  type slv83_vector  is array (natural range<>) of std_logic_vector( 82 downto 0);
  type slv84_vector  is array (natural range<>) of std_logic_vector( 83 downto 0);
  type slv85_vector  is array (natural range<>) of std_logic_vector( 84 downto 0);
  type slv86_vector  is array (natural range<>) of std_logic_vector( 85 downto 0);
  type slv87_vector  is array (natural range<>) of std_logic_vector( 86 downto 0);
  type slv88_vector  is array (natural range<>) of std_logic_vector( 87 downto 0);
  type slv89_vector  is array (natural range<>) of std_logic_vector( 88 downto 0);
  type slv90_vector  is array (natural range<>) of std_logic_vector( 89 downto 0);
  type slv91_vector  is array (natural range<>) of std_logic_vector( 90 downto 0);
  type slv92_vector  is array (natural range<>) of std_logic_vector( 91 downto 0);
  type slv93_vector  is array (natural range<>) of std_logic_vector( 92 downto 0);
  type slv94_vector  is array (natural range<>) of std_logic_vector( 93 downto 0);
  type slv95_vector  is array (natural range<>) of std_logic_vector( 94 downto 0);
  type slv96_vector  is array (natural range<>) of std_logic_vector( 95 downto 0);
  type slv97_vector  is array (natural range<>) of std_logic_vector( 96 downto 0);
  type slv98_vector  is array (natural range<>) of std_logic_vector( 97 downto 0);
  type slv99_vector  is array (natural range<>) of std_logic_vector( 98 downto 0);
  type slv100_vector is array (natural range<>) of std_logic_vector( 99 downto 0);
  type slv101_vector is array (natural range<>) of std_logic_vector(100 downto 0);
  type slv102_vector is array (natural range<>) of std_logic_vector(101 downto 0);
  type slv103_vector is array (natural range<>) of std_logic_vector(102 downto 0);
  type slv104_vector is array (natural range<>) of std_logic_vector(103 downto 0);
  type slv105_vector is array (natural range<>) of std_logic_vector(104 downto 0);
  type slv106_vector is array (natural range<>) of std_logic_vector(105 downto 0);
  type slv107_vector is array (natural range<>) of std_logic_vector(106 downto 0);
  type slv108_vector is array (natural range<>) of std_logic_vector(107 downto 0);
  type slv109_vector is array (natural range<>) of std_logic_vector(108 downto 0);
  type slv110_vector is array (natural range<>) of std_logic_vector(109 downto 0);
  type slv111_vector is array (natural range<>) of std_logic_vector(110 downto 0);
  type slv112_vector is array (natural range<>) of std_logic_vector(111 downto 0);
  type slv113_vector is array (natural range<>) of std_logic_vector(112 downto 0);
  type slv114_vector is array (natural range<>) of std_logic_vector(113 downto 0);
  type slv115_vector is array (natural range<>) of std_logic_vector(114 downto 0);
  type slv116_vector is array (natural range<>) of std_logic_vector(115 downto 0);
  type slv117_vector is array (natural range<>) of std_logic_vector(116 downto 0);
  type slv118_vector is array (natural range<>) of std_logic_vector(117 downto 0);
  type slv119_vector is array (natural range<>) of std_logic_vector(118 downto 0);
  type slv120_vector is array (natural range<>) of std_logic_vector(119 downto 0);
  type slv121_vector is array (natural range<>) of std_logic_vector(120 downto 0);
  type slv122_vector is array (natural range<>) of std_logic_vector(121 downto 0);
  type slv123_vector is array (natural range<>) of std_logic_vector(122 downto 0);
  type slv124_vector is array (natural range<>) of std_logic_vector(123 downto 0);
  type slv125_vector is array (natural range<>) of std_logic_vector(124 downto 0);
  type slv126_vector is array (natural range<>) of std_logic_vector(125 downto 0);
  type slv127_vector is array (natural range<>) of std_logic_vector(126 downto 0);
  type slv128_vector is array (natural range<>) of std_logic_vector(127 downto 0);
  type slv129_vector is array (natural range<>) of std_logic_vector(128 downto 0);
  type slv130_vector is array (natural range<>) of std_logic_vector(129 downto 0);
  type slv131_vector is array (natural range<>) of std_logic_vector(130 downto 0);
  type slv132_vector is array (natural range<>) of std_logic_vector(131 downto 0);
  type slv133_vector is array (natural range<>) of std_logic_vector(132 downto 0);
  type slv134_vector is array (natural range<>) of std_logic_vector(133 downto 0);
  type slv135_vector is array (natural range<>) of std_logic_vector(134 downto 0);
  type slv136_vector is array (natural range<>) of std_logic_vector(135 downto 0);
  type slv137_vector is array (natural range<>) of std_logic_vector(136 downto 0);
  type slv138_vector is array (natural range<>) of std_logic_vector(137 downto 0);
  type slv139_vector is array (natural range<>) of std_logic_vector(138 downto 0);
  type slv140_vector is array (natural range<>) of std_logic_vector(139 downto 0);
  type slv141_vector is array (natural range<>) of std_logic_vector(140 downto 0);
  type slv142_vector is array (natural range<>) of std_logic_vector(141 downto 0);
  type slv143_vector is array (natural range<>) of std_logic_vector(142 downto 0);
  type slv144_vector is array (natural range<>) of std_logic_vector(143 downto 0);
  type slv145_vector is array (natural range<>) of std_logic_vector(144 downto 0);
  type slv146_vector is array (natural range<>) of std_logic_vector(145 downto 0);
  type slv147_vector is array (natural range<>) of std_logic_vector(146 downto 0);
  type slv148_vector is array (natural range<>) of std_logic_vector(147 downto 0);
  type slv149_vector is array (natural range<>) of std_logic_vector(148 downto 0);
  type slv150_vector is array (natural range<>) of std_logic_vector(149 downto 0);
  type slv151_vector is array (natural range<>) of std_logic_vector(150 downto 0);
  type slv152_vector is array (natural range<>) of std_logic_vector(151 downto 0);
  type slv153_vector is array (natural range<>) of std_logic_vector(152 downto 0);
  type slv154_vector is array (natural range<>) of std_logic_vector(153 downto 0);
  type slv155_vector is array (natural range<>) of std_logic_vector(154 downto 0);
  type slv156_vector is array (natural range<>) of std_logic_vector(155 downto 0);
  type slv157_vector is array (natural range<>) of std_logic_vector(156 downto 0);
  type slv158_vector is array (natural range<>) of std_logic_vector(157 downto 0);
  type slv159_vector is array (natural range<>) of std_logic_vector(158 downto 0);
  type slv160_vector is array (natural range<>) of std_logic_vector(159 downto 0);
  type slv161_vector is array (natural range<>) of std_logic_vector(160 downto 0);
  type slv162_vector is array (natural range<>) of std_logic_vector(161 downto 0);
  type slv163_vector is array (natural range<>) of std_logic_vector(162 downto 0);
  type slv164_vector is array (natural range<>) of std_logic_vector(163 downto 0);
  type slv165_vector is array (natural range<>) of std_logic_vector(164 downto 0);
  type slv166_vector is array (natural range<>) of std_logic_vector(165 downto 0);
  type slv167_vector is array (natural range<>) of std_logic_vector(166 downto 0);
  type slv168_vector is array (natural range<>) of std_logic_vector(167 downto 0);
  type slv169_vector is array (natural range<>) of std_logic_vector(168 downto 0);
  type slv170_vector is array (natural range<>) of std_logic_vector(169 downto 0);
  type slv171_vector is array (natural range<>) of std_logic_vector(170 downto 0);
  type slv172_vector is array (natural range<>) of std_logic_vector(171 downto 0);
  type slv173_vector is array (natural range<>) of std_logic_vector(172 downto 0);
  type slv174_vector is array (natural range<>) of std_logic_vector(173 downto 0);
  type slv175_vector is array (natural range<>) of std_logic_vector(174 downto 0);
  type slv176_vector is array (natural range<>) of std_logic_vector(175 downto 0);
  type slv177_vector is array (natural range<>) of std_logic_vector(176 downto 0);
  type slv178_vector is array (natural range<>) of std_logic_vector(177 downto 0);
  type slv179_vector is array (natural range<>) of std_logic_vector(178 downto 0);
  type slv180_vector is array (natural range<>) of std_logic_vector(179 downto 0);
  type slv181_vector is array (natural range<>) of std_logic_vector(180 downto 0);
  type slv182_vector is array (natural range<>) of std_logic_vector(181 downto 0);
  type slv183_vector is array (natural range<>) of std_logic_vector(182 downto 0);
  type slv184_vector is array (natural range<>) of std_logic_vector(183 downto 0);
  type slv185_vector is array (natural range<>) of std_logic_vector(184 downto 0);
  type slv186_vector is array (natural range<>) of std_logic_vector(185 downto 0);
  type slv187_vector is array (natural range<>) of std_logic_vector(186 downto 0);
  type slv188_vector is array (natural range<>) of std_logic_vector(187 downto 0);
  type slv189_vector is array (natural range<>) of std_logic_vector(188 downto 0);
  type slv190_vector is array (natural range<>) of std_logic_vector(189 downto 0);
  type slv191_vector is array (natural range<>) of std_logic_vector(190 downto 0);
  type slv192_vector is array (natural range<>) of std_logic_vector(191 downto 0);
  type slv193_vector is array (natural range<>) of std_logic_vector(192 downto 0);
  type slv194_vector is array (natural range<>) of std_logic_vector(193 downto 0);
  type slv195_vector is array (natural range<>) of std_logic_vector(194 downto 0);
  type slv196_vector is array (natural range<>) of std_logic_vector(195 downto 0);
  type slv197_vector is array (natural range<>) of std_logic_vector(196 downto 0);
  type slv198_vector is array (natural range<>) of std_logic_vector(197 downto 0);
  type slv199_vector is array (natural range<>) of std_logic_vector(198 downto 0);
  type slv200_vector is array (natural range<>) of std_logic_vector(199 downto 0);
  type slv201_vector is array (natural range<>) of std_logic_vector(200 downto 0);
  type slv202_vector is array (natural range<>) of std_logic_vector(201 downto 0);
  type slv203_vector is array (natural range<>) of std_logic_vector(202 downto 0);
  type slv204_vector is array (natural range<>) of std_logic_vector(203 downto 0);
  type slv205_vector is array (natural range<>) of std_logic_vector(204 downto 0);
  type slv206_vector is array (natural range<>) of std_logic_vector(205 downto 0);
  type slv207_vector is array (natural range<>) of std_logic_vector(206 downto 0);
  type slv208_vector is array (natural range<>) of std_logic_vector(207 downto 0);
  type slv209_vector is array (natural range<>) of std_logic_vector(208 downto 0);
  type slv210_vector is array (natural range<>) of std_logic_vector(209 downto 0);
  type slv211_vector is array (natural range<>) of std_logic_vector(210 downto 0);
  type slv212_vector is array (natural range<>) of std_logic_vector(211 downto 0);
  type slv213_vector is array (natural range<>) of std_logic_vector(212 downto 0);
  type slv214_vector is array (natural range<>) of std_logic_vector(213 downto 0);
  type slv215_vector is array (natural range<>) of std_logic_vector(214 downto 0);
  type slv216_vector is array (natural range<>) of std_logic_vector(215 downto 0);
  type slv217_vector is array (natural range<>) of std_logic_vector(216 downto 0);
  type slv218_vector is array (natural range<>) of std_logic_vector(217 downto 0);
  type slv219_vector is array (natural range<>) of std_logic_vector(218 downto 0);
  type slv220_vector is array (natural range<>) of std_logic_vector(219 downto 0);
  type slv221_vector is array (natural range<>) of std_logic_vector(220 downto 0);
  type slv222_vector is array (natural range<>) of std_logic_vector(221 downto 0);
  type slv223_vector is array (natural range<>) of std_logic_vector(222 downto 0);
  type slv224_vector is array (natural range<>) of std_logic_vector(223 downto 0);
  type slv225_vector is array (natural range<>) of std_logic_vector(224 downto 0);
  type slv226_vector is array (natural range<>) of std_logic_vector(225 downto 0);
  type slv227_vector is array (natural range<>) of std_logic_vector(226 downto 0);
  type slv228_vector is array (natural range<>) of std_logic_vector(227 downto 0);
  type slv229_vector is array (natural range<>) of std_logic_vector(228 downto 0);
  type slv230_vector is array (natural range<>) of std_logic_vector(229 downto 0);
  type slv231_vector is array (natural range<>) of std_logic_vector(230 downto 0);
  type slv232_vector is array (natural range<>) of std_logic_vector(231 downto 0);
  type slv233_vector is array (natural range<>) of std_logic_vector(232 downto 0);
  type slv234_vector is array (natural range<>) of std_logic_vector(233 downto 0);
  type slv235_vector is array (natural range<>) of std_logic_vector(234 downto 0);
  type slv236_vector is array (natural range<>) of std_logic_vector(235 downto 0);
  type slv237_vector is array (natural range<>) of std_logic_vector(236 downto 0);
  type slv238_vector is array (natural range<>) of std_logic_vector(237 downto 0);
  type slv239_vector is array (natural range<>) of std_logic_vector(238 downto 0);
  type slv240_vector is array (natural range<>) of std_logic_vector(239 downto 0);
  type slv241_vector is array (natural range<>) of std_logic_vector(240 downto 0);
  type slv242_vector is array (natural range<>) of std_logic_vector(241 downto 0);
  type slv243_vector is array (natural range<>) of std_logic_vector(242 downto 0);
  type slv244_vector is array (natural range<>) of std_logic_vector(243 downto 0);
  type slv245_vector is array (natural range<>) of std_logic_vector(244 downto 0);
  type slv246_vector is array (natural range<>) of std_logic_vector(245 downto 0);
  type slv247_vector is array (natural range<>) of std_logic_vector(246 downto 0);
  type slv248_vector is array (natural range<>) of std_logic_vector(247 downto 0);
  type slv249_vector is array (natural range<>) of std_logic_vector(248 downto 0);
  type slv250_vector is array (natural range<>) of std_logic_vector(249 downto 0);
  type slv251_vector is array (natural range<>) of std_logic_vector(250 downto 0);
  type slv252_vector is array (natural range<>) of std_logic_vector(251 downto 0);
  type slv253_vector is array (natural range<>) of std_logic_vector(252 downto 0);
  type slv254_vector is array (natural range<>) of std_logic_vector(253 downto 0);
  type slv255_vector is array (natural range<>) of std_logic_vector(254 downto 0);
  type slv256_vector is array (natural range<>) of std_logic_vector(255 downto 0);

  type int_vector    is array (natural range<>) of integer;

  type bool_vector   is array (natural range<>) of boolean;

  subtype uint1  is integer range 0 to          1;
  subtype uint2  is integer range 0 to          3;
  subtype uint3  is integer range 0 to          7;
  subtype uint4  is integer range 0 to         15;
  subtype uint5  is integer range 0 to         31;
  subtype uint6  is integer range 0 to         63;
  subtype uint7  is integer range 0 to        127;
  subtype uint8  is integer range 0 to        255;
  subtype uint9  is integer range 0 to        511;
  subtype uint10 is integer range 0 to       1023;
  subtype uint11 is integer range 0 to       2047;
  subtype uint12 is integer range 0 to       4095;
  subtype uint13 is integer range 0 to       8191;
  subtype uint14 is integer range 0 to      16383;
  subtype uint15 is integer range 0 to      32767;
  subtype uint16 is integer range 0 to      65535;
  subtype uint17 is integer range 0 to     131071;
  subtype uint18 is integer range 0 to     262143;
  subtype uint19 is integer range 0 to     524287;
  subtype uint20 is integer range 0 to    1048575;
  subtype uint21 is integer range 0 to    2097151;
  subtype uint22 is integer range 0 to    4194303;
  subtype uint23 is integer range 0 to    8388607;
  subtype uint24 is integer range 0 to   16777215;
  subtype uint25 is integer range 0 to   33554431;
  subtype uint26 is integer range 0 to   67108863;
  subtype uint27 is integer range 0 to  134217727;
  subtype uint28 is integer range 0 to  268435455;
  subtype uint29 is integer range 0 to  536870911;
  subtype uint30 is integer range 0 to 1073741823;
  subtype uint31 is integer range 0 to 2147483647;

  subtype sint2  is integer range          -2 to          1;
  subtype sint3  is integer range          -4 to          3;
  subtype sint4  is integer range          -8 to          7;
  subtype sint5  is integer range         -16 to         15;
  subtype sint6  is integer range         -32 to         31;
  subtype sint7  is integer range         -64 to         63;
  subtype sint8  is integer range        -128 to        127;
  subtype sint9  is integer range        -256 to        255;
  subtype sint10 is integer range        -512 to        511;
  subtype sint11 is integer range       -1024 to       1023;
  subtype sint12 is integer range       -2048 to       2047;
  subtype sint13 is integer range       -4096 to       4095;
  subtype sint14 is integer range       -8192 to       8191;
  subtype sint15 is integer range      -16384 to      16383;
  subtype sint16 is integer range      -32768 to      32767;
  subtype sint17 is integer range      -65536 to      65535;
  subtype sint18 is integer range     -131072 to     131071;
  subtype sint19 is integer range     -262144 to     262143;
  subtype sint20 is integer range     -524288 to     524287;
  subtype sint21 is integer range    -1048576 to    1048575;
  subtype sint22 is integer range    -2097152 to    2097151;
  subtype sint23 is integer range    -4194304 to    4194303;
  subtype sint24 is integer range    -8388608 to    8388607;
  subtype sint25 is integer range   -16777216 to   16777215;
  subtype sint26 is integer range   -33554432 to   33554431;
  subtype sint27 is integer range   -67108864 to   67108863;
  subtype sint28 is integer range  -134217728 to  134217727;
  subtype sint29 is integer range  -268435456 to  268435455;
  subtype sint30 is integer range  -536870912 to  536870911;
  subtype sint31 is integer range -1073741824 to 1073741823;
end typ;
